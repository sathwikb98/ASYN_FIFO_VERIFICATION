`define DSIZE 8 // size of data bus
`define ASIZE 4 // size of address bus
`define no_of_transaction 10
