`define DSIZE 8 // size of data bus
`define ASIZE 4 // size of address
`define DEPTH 16  // depth of fifo memory !
`define no_of_transaction 50
