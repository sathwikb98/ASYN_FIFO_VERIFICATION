package asyn_fifo_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "defines.svh"

  `include "fifo_write_seq_item.sv" // sequence item !
  `include "fifo_read_seq_item.sv"

  `include "fifo_write_sequence.sv" // sequence 
  `include "fifo_read_sequence.sv"
  
  `include "fifo_write_sequencer.sv" // sequencer 
  `include "fifo_read_sequencer.sv"

  `include "fifo_write_driver.sv" // driver  !
  `include "fifo_read_driver.sv"

  `include "fifo_write_monitor.sv" // monitor !
  `include "fifo_read_monitor.sv"

  `include "fifo_scoreboard.sv" 
  `include "fifo_subscriber.sv"

  `include "fifo_write_agent.sv"
  `include "fifo_read_agent.sv"

  `include "fifo_virtual_sequencer.sv"
  
  `include "fifo_env.sv"
  
  `include "fifo_virtual_sequence.sv" // virtual sequencer !
  
  `include "fifo_test.sv"
  
endpackage
